LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

entity LUT_encoder is
port (
    F	:	in STD_LOGIC_VECTOR(127 downto 0);
    s	: 	out STD_LOGIC_VECTOR(7 downto 0)
    );
end LUT_encoder;	

architecture tabla of LUT_encoder is
	begin
		process(F)
		begin case F is
		
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001" => s <= "00000000";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010" => s <= "00000001";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100" => s <= "00000010";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000" => s <= "00000011";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000" => s <= "00000100";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000" => s <= "00000101";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000" => s <= "00000110";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000" => s <= "00000111";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000" => s <= "00001000";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000" => s <= "00001001";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000" => s <= "00001010";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000" => s <= "00001011";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000" => s <= "00001100";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000" => s <= "00001101";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000" => s <= "00001110";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000" => s <= "00001111";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000" => s <= "00010000";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000" => s <= "00010001";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000" => s <= "00010010";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000" => s <= "00010011";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000" => s <= "00010100";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000" => s <= "00010101";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000" => s <= "00010110";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000" => s <= "00010111";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000" => s <= "00011000";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000" => s <= "00011001";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000" => s <= "00011010";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000" => s <= "00011011";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000" => s <= "00011100";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000" => s <= "00011101";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000" => s <= "00011110";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000" => s <= "00011111";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000" => s <= "00100000";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000" => s <= "00100001";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000" => s <= "00100010";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000" => s <= "00100011";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000" => s <= "00100100";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000" => s <= "00100101";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000" => s <= "00100110";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000" => s <= "00100111";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000" => s <= "00101000";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000" => s <= "00101001";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000" => s <= "00101010";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000" => s <= "00101011";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000" => s <= "00101100";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000" => s <= "00101101";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000" => s <= "00101110";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000" => s <= "00101111";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000" => s <= "00110000";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000" => s <= "00110001";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000" => s <= "00110010";
when "00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000" => s <= "00110011";
when "00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000" => s <= "00110100";
when "00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000" => s <= "00110101";
when "00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000" => s <= "00110110";
when "00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000" => s <= "00110111";
when "00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000" => s <= "00111000";
when "00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000" => s <= "00111001";
when "00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000" => s <= "00111010";
when "00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000" => s <= "00111011";
when "00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000" => s <= "00111100";
when "00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000" => s <= "00111101";
when "00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000" => s <= "00111110";
when "00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000" => s <= "00111111";
when "00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000" => s <= "01000000";
when "00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000" => s <= "01000001";
when "00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000" => s <= "01000010";
when "00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000" => s <= "01000011";
when "00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000" => s <= "01000100";
when "00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01000101";
when "00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01000110";
when "00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01000111";
when "00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01001000";
when "00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01001001";
when "00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01001010";
when "00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01001011";
when "00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01001100";
when "00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01001101";
when "00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01001110";
when "00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01001111";
when "00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01010000";
when "00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01010001";
when "00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01010010";
when "00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01010011";
when "00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01010100";
when "00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01010101";
when "00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01010110";
when "00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01010111";
when "00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01011000";
when "00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01011001";
when "00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01011010";
when "00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01011011";
when "00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01011100";
when "00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01011101";
when "00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01011110";
when "00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01011111";
when "00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01100000";
when "00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01100001";
when "00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01100010";
when "00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01100011";
when "00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01100100";
when "00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01100101";
when "00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01100110";
when "00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01100111";
when "00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01101000";
when "00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01101001";
when "00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01101010";
when "00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01101011";
when "00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01101100";
when "00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01101101";
when "00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01101110";
when "00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01101111";
when "00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01110000";
when "00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01110001";
when "00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01110010";
when "00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01110011";
when "00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01110100";
when "00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01110101";
when "00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01110110";
when "00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01110111";
when "00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01111000";
when "00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01111001";
when "00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01111010";
when "00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01111011";
when "00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01111100";
when "00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01111101";
when "01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01111110";
when "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "01111111";
when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" => s <= "10000000";	  
when others => s <="11111111";
      end case;
   end process;
end tabla;